LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.ALL;

PACKAGE MIPS_Types IS
	SUBTYPE BYTE IS STD_LOGIC_VECTOR (7 DOWNTO 0);
	SUBTYPE WORD IS STD_LOGIC_VECTOR (15 DOWNTO 0);
	SUBTYPE REG_ADDRESS IS STD_LOGIC_VECTOR (2 DOWNTO 0);
	
	TYPE ALU_OP IS (AND_OP, ADD_OP, ADDU_OP, SUB_OP, CAS_OP, SHL_OP, SHR_OP, UNDEFINED);
	TYPE INST_OP IS (ZERO, ANDI, ADDI, SLTI, LW, LLB, SW, SLB, LWS, BEQ, BNE,
	J, JAL, JALR, LUI, TERMINATE);
	TYPE MEM_INST IS ARRAY (0 TO 2**16 - 1) OF WORD;
	TYPE MEM_DATA IS ARRAY (0 TO 2**16 - 1)	OF BYTE;
	TYPE REG_FILE IS ARRAY (0 TO 7) OF WORD;
	
	TYPE RTYPE_INSTRUCTION IS RECORD
		OPCODE : INST_OP;
		Rs: REG_ADDRESS;
		Rt: REG_ADDRESS;
		Rd: REG_ADDRESS;
		FUNC: STD_LOGIC_VECTOR (2 DOWNTO 0);
	END RECORD;
	
	TYPE ITYPE_INSTRUCTION IS RECORD
		OPCODE : INST_OP;
		Rs: REG_ADDRESS;
		Rt: REG_ADDRESS;
		Immediate: STD_LOGIC_VECTOR (5 DOWNTO 0);
	END RECORD;
	
	TYPE JTYPE_INSTRUCTION IS RECORD
		OPCODE : INST_OP;
		Immediate: STD_LOGIC_VECTOR (11 DOWNTO 0);
	END RECORD;
	
	FUNCTION MAX(a, b: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;
	FUNCTION RConv(Instruction: WORD) RETURN RTYPE_INSTRUCTION;
	FUNCTION IConv(Instruction: WORD) RETURN ITYPE_INSTRUCTION;
	FUNCTION JConv(Instruction: WORD) RETURN JTYPE_INSTRUCTION;
END PACKAGE MIPS_Types;

PACKAGE BODY MIPS_Types IS
	FUNCTION MAX(a, b: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
	BEGIN
		IF a > b THEN
			RETURN a;
		ELSE
			RETURN b;
		END IF;
	END FUNCTION MAX;
	
	FUNCTION RConv(Instruction: WORD) RETURN RTYPE_INSTRUCTION IS
	VARIABLE RInst: RTYPE_INSTRUCTION;
	BEGIN
		RInst.OPCODE := INST_OP'VAL(conv_integer(Instruction(15 DOWNTO 12)));
		RInst.Rs := Instruction(11 DOWNTO 9);
		RInst.Rt := Instruction(8 DOWNTO 6);
		RInst.Rd := Instruction(5 DOWNTO 3);
		RInst.FUNC := Instruction(2 DOWNTO 0);
		RETURN RInst;
	END FUNCTION RConv;
	
	FUNCTION IConv(Instruction: WORD) RETURN ITYPE_INSTRUCTION IS
	VARIABLE IInst: ITYPE_INSTRUCTION;
	BEGIN
		IInst.OPCODE := INST_OP'VAL(conv_integer(Instruction(15 DOWNTO 12)));
		IInst.Rs := Instruction(11 DOWNTO 9);
		IInst.Rt := Instruction(8 DOWNTO 6);
		IInst.Immediate := Instruction(5 DOWNTO 0);
		RETURN IInst;
	END FUNCTION IConv;
	
	FUNCTION JConv(Instruction: WORD) RETURN JTYPE_INSTRUCTION IS
	VARIABLE JInst: JTYPE_INSTRUCTION;
	BEGIN
		JInst.OPCODE := INST_OP'VAL(conv_integer(Instruction(15 DOWNTO 12)));
		JInst.Immediate := Instruction(11 DOWNTO 0);
		RETURN JInst;
	END FUNCTION JConv;
	
END PACKAGE BODY MIPS_Types;